module setbit (A);
  output A;
  wire A;

  assign A = 1;

endmodule
